magic
tech sky130A
magscale 1 2
timestamp 1692670061
<< error_s >>
rect 129 1029 187 1035
rect 129 995 141 1029
rect 129 989 187 995
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect -28 -28 -21 100
rect 0 0 7 128
rect -29 -138 29 -132
rect -29 -172 -17 -138
rect -29 -178 29 -172
rect 0 -206 57 -200
<< pwell >>
rect -211 -310 211 310
<< nmos >>
rect -15 -100 15 100
<< ndiff >>
rect -73 88 -15 100
rect -73 -88 -61 88
rect -27 -88 -15 88
rect -73 -100 -15 -88
rect 15 88 73 100
rect 15 -88 27 88
rect 61 -88 73 88
rect 15 -100 73 -88
<< ndiffc >>
rect -61 -88 -27 88
rect 27 -88 61 88
<< psubdiff >>
rect -175 240 -79 274
rect 79 240 175 274
rect -175 178 -141 240
rect 141 178 175 240
rect -175 -240 -141 -178
rect 141 -240 175 -178
rect -175 -274 -79 -240
rect 79 -274 175 -240
<< psubdiffcont >>
rect -79 240 79 274
rect -175 -178 -141 178
rect 141 -178 175 178
rect -79 -274 79 -240
<< poly >>
rect -33 172 33 188
rect -33 138 -17 172
rect 17 138 33 172
rect -33 122 33 138
rect -15 100 15 122
rect -15 -122 15 -100
rect -33 -138 33 -122
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect -33 -188 33 -172
<< polycont >>
rect -17 138 17 172
rect -17 -172 17 -138
<< locali >>
rect -175 240 -79 274
rect 79 240 175 274
rect -175 178 -141 240
rect 141 178 175 240
rect -33 138 -17 172
rect 17 138 33 172
rect -61 88 -27 104
rect -61 -104 -27 -88
rect 27 88 61 104
rect 27 -104 61 -88
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect -175 -240 -141 -178
rect 141 -240 175 -178
rect -175 -274 -79 -240
rect 79 -274 175 -240
<< viali >>
rect -17 138 17 172
rect -175 -120 -141 120
rect -61 -88 -27 88
rect 27 -88 61 88
rect -17 -172 17 -138
<< metal1 >>
rect 0 178 200 200
rect -29 172 200 178
rect -29 138 -17 172
rect 17 138 200 172
rect -29 132 200 138
rect -181 120 -135 132
rect -181 -120 -175 120
rect -141 -120 -135 120
rect -67 88 -21 100
rect -67 -88 -61 88
rect -27 -88 -21 88
rect 0 88 200 132
rect 0 0 27 88
rect -67 -100 -21 -88
rect 21 -88 27 0
rect 61 0 200 88
rect 61 -88 67 0
rect 21 -100 67 -88
rect -181 -132 -135 -120
rect -29 -138 29 -132
rect -29 -172 -17 -138
rect 17 -172 29 -138
rect -29 -178 29 -172
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__nfet_01v8_648S5X  X0
timestamp 1692470706
transform 1 0 158 0 1 857
box -211 -310 211 310
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 a_n73_n100#
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 a_n33_n188#
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 a_15_n100#
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 a_n175_n274#
port 3 nsew
<< properties >>
string FIXED_BBOX -158 -257 158 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 50 viagt 0
<< end >>
